magic
tech sky130A
timestamp 1760114222
<< nmos >>
rect -40 70 -25 120
rect 10 70 25 140
rect 65 70 80 120
rect 125 70 140 140
rect -40 -180 -25 -130
rect 10 -180 25 -110
rect 65 -180 80 -130
rect 125 -180 140 -110
<< ndiff >>
rect -15 120 10 140
rect -85 105 -40 120
rect -85 85 -70 105
rect -50 85 -40 105
rect -85 70 -40 85
rect -25 70 10 120
rect 25 120 55 140
rect 100 120 125 140
rect 25 105 65 120
rect 25 85 35 105
rect 55 85 65 105
rect 25 70 65 85
rect 80 105 125 120
rect 80 85 95 105
rect 115 85 125 105
rect 80 70 125 85
rect 140 70 165 140
rect -15 -130 10 -110
rect -85 -145 -40 -130
rect -85 -165 -70 -145
rect -50 -165 -40 -145
rect -85 -180 -40 -165
rect -25 -180 10 -130
rect 25 -130 55 -110
rect 100 -130 125 -110
rect 25 -145 65 -130
rect 25 -165 35 -145
rect 55 -165 65 -145
rect 25 -180 65 -165
rect 80 -145 125 -130
rect 80 -165 95 -145
rect 115 -165 125 -145
rect 80 -180 125 -165
rect 140 -180 165 -110
<< ndiffc >>
rect -70 85 -50 105
rect 35 85 55 105
rect 95 85 115 105
rect -70 -165 -50 -145
rect 35 -165 55 -145
rect 95 -165 115 -145
<< psubdiff >>
rect -135 105 -85 120
rect -135 85 -120 105
rect -100 85 -85 105
rect -135 70 -85 85
rect -135 -145 -85 -130
rect -135 -165 -120 -145
rect -100 -165 -85 -145
rect -135 -180 -85 -165
<< psubdiffcont >>
rect -120 85 -100 105
rect -120 -165 -100 -145
<< poly >>
rect 10 140 25 155
rect -40 120 -25 135
rect 65 120 80 155
rect 125 140 140 155
rect -40 -130 -25 70
rect 10 55 25 70
rect 0 10 40 55
rect 0 -95 40 -50
rect 10 -110 25 -95
rect 65 -130 80 70
rect 125 55 140 70
rect 125 -110 140 -95
rect -40 -195 -25 -180
rect 10 -195 25 -180
rect 65 -195 80 -180
rect 125 -195 140 -180
<< locali >>
rect -130 105 -40 115
rect -130 85 -120 105
rect -100 85 -70 105
rect -50 85 -40 105
rect -130 75 -40 85
rect 25 105 65 115
rect 25 85 35 105
rect 55 85 65 105
rect 25 75 65 85
rect 85 105 125 115
rect 85 85 95 105
rect 115 85 125 105
rect 85 75 125 85
rect -130 -145 -40 -135
rect -130 -165 -120 -145
rect -100 -165 -70 -145
rect -50 -165 -40 -145
rect -130 -175 -40 -165
rect 25 -145 65 -135
rect 25 -165 35 -145
rect 55 -165 65 -145
rect 25 -175 65 -165
rect 85 -145 125 -135
rect 85 -165 95 -145
rect 115 -165 125 -145
rect 85 -175 125 -165
<< end >>
