magic
tech sky130A
timestamp 1760147834
<< nwell >>
rect 90 530 180 610
rect -95 70 330 530
<< nmos >>
rect -10 -55 5 -5
rect 50 -55 65 -5
rect 160 -110 175 -5
rect 270 -55 285 -5
rect -10 -315 5 -265
rect 50 -315 65 -265
rect 160 -315 175 -205
rect 270 -315 285 -265
<< pmos >>
rect -10 405 5 510
rect 90 405 105 510
rect 160 405 175 510
rect 225 405 240 510
rect -10 90 5 195
rect 90 90 105 195
rect 160 90 175 195
rect 225 90 240 195
<< ndiff >>
rect -60 -20 -10 -5
rect -60 -40 -45 -20
rect -25 -40 -10 -20
rect -60 -55 -10 -40
rect 5 -20 50 -5
rect 5 -40 15 -20
rect 35 -40 50 -20
rect 5 -55 50 -40
rect 65 -20 160 -5
rect 65 -40 85 -20
rect 140 -40 160 -20
rect 65 -55 160 -40
rect 135 -110 160 -55
rect 175 -20 270 -5
rect 175 -40 200 -20
rect 255 -40 270 -20
rect 175 -55 270 -40
rect 285 -20 330 -5
rect 285 -40 300 -20
rect 320 -40 330 -20
rect 285 -55 330 -40
rect 175 -110 200 -55
rect 135 -265 160 -205
rect -60 -280 -10 -265
rect -60 -300 -45 -280
rect -25 -300 -10 -280
rect -60 -315 -10 -300
rect 5 -280 50 -265
rect 5 -300 15 -280
rect 35 -300 50 -280
rect 5 -315 50 -300
rect 65 -280 160 -265
rect 65 -300 85 -280
rect 140 -300 160 -280
rect 65 -315 160 -300
rect 175 -265 200 -205
rect 175 -280 270 -265
rect 175 -300 200 -280
rect 255 -300 270 -280
rect 175 -315 270 -300
rect 285 -280 330 -265
rect 285 -300 300 -280
rect 320 -300 330 -280
rect 285 -315 330 -300
<< pdiff >>
rect -60 495 -10 510
rect -60 420 -40 495
rect -20 420 -10 495
rect -60 405 -10 420
rect 5 495 90 510
rect 5 420 60 495
rect 80 420 90 495
rect 5 405 90 420
rect 105 495 160 510
rect 105 420 130 495
rect 150 420 160 495
rect 105 405 160 420
rect 175 495 225 510
rect 175 420 190 495
rect 210 420 225 495
rect 175 405 225 420
rect 240 495 285 510
rect 240 420 250 495
rect 270 420 285 495
rect 240 405 285 420
rect -60 180 -10 195
rect -60 105 -40 180
rect -20 105 -10 180
rect -60 90 -10 105
rect 5 180 90 195
rect 5 105 60 180
rect 80 105 90 180
rect 5 90 90 105
rect 105 180 160 195
rect 105 105 130 180
rect 150 105 160 180
rect 105 90 160 105
rect 175 180 225 195
rect 175 105 190 180
rect 210 105 225 180
rect 175 90 225 105
rect 240 180 285 195
rect 240 105 250 180
rect 270 105 285 180
rect 240 90 285 105
<< ndiffc >>
rect -45 -40 -25 -20
rect 15 -40 35 -20
rect 85 -40 140 -20
rect 200 -40 255 -20
rect 300 -40 320 -20
rect -45 -300 -25 -280
rect 15 -300 35 -280
rect 85 -300 140 -280
rect 200 -300 255 -280
rect 300 -300 320 -280
<< pdiffc >>
rect -40 420 -20 495
rect 60 420 80 495
rect 130 420 150 495
rect 190 420 210 495
rect 250 420 270 495
rect -40 105 -20 180
rect 60 105 80 180
rect 130 105 150 180
rect 190 105 210 180
rect 250 105 270 180
<< psubdiff >>
rect -70 -140 -20 -125
rect -70 -160 -55 -140
rect -35 -160 -20 -140
rect -70 -175 -20 -160
<< nsubdiff >>
rect 110 575 160 590
rect 110 555 125 575
rect 145 555 160 575
rect 110 540 160 555
<< psubdiffcont >>
rect -55 -160 -35 -140
<< nsubdiffcont >>
rect 125 555 145 575
<< poly >>
rect -10 510 5 525
rect 90 510 105 525
rect 160 510 175 525
rect 225 510 240 525
rect -10 195 5 405
rect 90 395 105 405
rect 30 380 105 395
rect 30 285 45 380
rect 70 340 125 350
rect 70 320 80 340
rect 100 320 125 340
rect 70 310 125 320
rect 30 275 85 285
rect 30 255 55 275
rect 75 255 85 275
rect 30 245 85 255
rect 110 220 125 310
rect 90 205 125 220
rect 90 195 105 205
rect 160 195 175 405
rect 225 395 240 405
rect 225 380 300 395
rect 205 340 260 350
rect 205 320 230 340
rect 250 320 260 340
rect 205 310 260 320
rect 205 220 220 310
rect 285 285 300 380
rect 245 275 300 285
rect 245 255 255 275
rect 275 255 300 275
rect 245 245 300 255
rect 205 205 240 220
rect 225 195 240 205
rect -10 60 5 90
rect -35 50 5 60
rect -35 30 -25 50
rect -5 30 5 50
rect 90 35 105 90
rect 160 60 175 90
rect -35 20 5 30
rect -10 -5 5 20
rect 50 20 105 35
rect 135 50 175 60
rect 135 30 145 50
rect 165 30 175 50
rect 135 20 175 30
rect 225 35 240 90
rect 225 20 285 35
rect 50 -5 65 20
rect 160 -5 175 20
rect 270 -5 285 20
rect -10 -265 5 -55
rect 50 -65 65 -55
rect 50 -80 125 -65
rect 30 -120 85 -110
rect 30 -140 55 -120
rect 75 -140 85 -120
rect 30 -150 85 -140
rect 30 -240 45 -150
rect 110 -175 125 -80
rect 270 -65 285 -55
rect 210 -80 285 -65
rect 70 -185 125 -175
rect 70 -205 80 -185
rect 100 -205 125 -185
rect 160 -205 175 -110
rect 210 -175 225 -80
rect 250 -120 305 -110
rect 250 -140 260 -120
rect 280 -140 305 -120
rect 250 -150 305 -140
rect 210 -185 265 -175
rect 210 -205 235 -185
rect 255 -205 265 -185
rect 70 -215 125 -205
rect 30 -255 65 -240
rect 50 -265 65 -255
rect 210 -215 265 -205
rect 290 -240 305 -150
rect 270 -255 305 -240
rect 270 -265 285 -255
rect -10 -330 5 -315
rect 50 -330 65 -315
rect 160 -330 175 -315
rect 270 -330 285 -315
<< polycont >>
rect 80 320 100 340
rect 55 255 75 275
rect 230 320 250 340
rect 255 255 275 275
rect -25 30 -5 50
rect 145 30 165 50
rect 55 -140 75 -120
rect 80 -205 100 -185
rect 260 -140 280 -120
rect 235 -205 255 -185
<< locali >>
rect 115 575 155 585
rect 115 555 125 575
rect 145 555 155 575
rect 115 545 155 555
rect -95 505 -75 525
rect 135 510 155 545
rect -95 495 -10 505
rect -95 485 -40 495
rect -50 420 -40 485
rect -20 420 -10 495
rect -50 410 -10 420
rect 50 495 90 505
rect 50 420 60 495
rect 80 420 90 495
rect 50 410 90 420
rect 120 495 160 510
rect 310 505 330 525
rect 120 420 130 495
rect 150 420 160 495
rect 120 410 160 420
rect 70 350 90 410
rect 70 340 110 350
rect 70 320 80 340
rect 100 320 110 340
rect 70 310 110 320
rect 45 275 85 285
rect 45 255 55 275
rect 75 255 85 275
rect 45 245 85 255
rect 65 190 85 245
rect 135 190 160 410
rect -95 180 -10 190
rect -95 170 -40 180
rect -50 105 -40 170
rect -20 105 -10 180
rect -50 95 -10 105
rect 50 180 90 190
rect 50 105 60 180
rect 80 105 90 180
rect 50 95 90 105
rect 120 180 160 190
rect 120 105 130 180
rect 150 105 160 180
rect 120 95 160 105
rect 180 495 220 505
rect 180 420 190 495
rect 210 420 220 495
rect 180 410 220 420
rect 240 495 330 505
rect 240 420 250 495
rect 270 480 330 495
rect 270 420 280 480
rect 240 410 280 420
rect 180 190 200 410
rect 240 350 260 410
rect 220 340 260 350
rect 220 320 230 340
rect 250 320 260 340
rect 220 310 260 320
rect 245 275 285 285
rect 245 255 255 275
rect 275 255 285 275
rect 245 245 285 255
rect 245 190 265 245
rect 180 180 220 190
rect 180 105 190 180
rect 210 105 220 180
rect 180 95 220 105
rect 240 180 330 190
rect 240 105 250 180
rect 270 165 330 180
rect 270 105 280 165
rect 240 95 280 105
rect -35 50 5 60
rect -35 30 -25 50
rect -5 30 5 50
rect -35 20 5 30
rect 65 -10 90 95
rect 135 50 175 60
rect 135 30 145 50
rect 165 30 175 50
rect 135 20 175 30
rect 240 -10 265 95
rect -55 -20 -15 -10
rect -55 -40 -45 -20
rect -25 -40 -15 -20
rect -55 -50 -15 -40
rect -35 -130 -15 -50
rect -65 -140 -15 -130
rect -65 -160 -55 -140
rect -35 -160 -15 -140
rect -65 -170 -15 -160
rect -35 -270 -15 -170
rect -55 -280 -15 -270
rect -55 -300 -45 -280
rect -25 -300 -15 -280
rect -55 -310 -15 -300
rect 5 -20 45 -10
rect 5 -40 15 -20
rect 35 -40 45 -20
rect 5 -50 45 -40
rect 65 -20 155 -10
rect 65 -40 85 -20
rect 140 -40 155 -20
rect 65 -50 155 -40
rect 180 -20 270 -10
rect 180 -40 200 -20
rect 255 -40 270 -20
rect 180 -50 270 -40
rect 290 -20 330 -10
rect 290 -40 300 -20
rect 320 -40 330 -20
rect 290 -50 330 -40
rect 5 -270 25 -50
rect 65 -110 85 -50
rect 45 -120 85 -110
rect 45 -140 55 -120
rect 75 -140 85 -120
rect 45 -150 85 -140
rect 250 -110 270 -50
rect 250 -120 290 -110
rect 250 -140 260 -120
rect 280 -140 290 -120
rect 250 -150 290 -140
rect 70 -185 110 -175
rect 70 -205 80 -185
rect 100 -205 110 -185
rect 70 -215 110 -205
rect 90 -270 110 -215
rect 225 -185 265 -175
rect 225 -205 235 -185
rect 255 -205 265 -185
rect 225 -215 265 -205
rect 225 -270 245 -215
rect 310 -270 330 -50
rect 5 -280 45 -270
rect 5 -300 15 -280
rect 35 -300 45 -280
rect 5 -310 45 -300
rect 65 -280 155 -270
rect 65 -300 85 -280
rect 140 -300 155 -280
rect 65 -310 155 -300
rect 180 -280 270 -270
rect 180 -300 200 -280
rect 255 -300 270 -280
rect 180 -310 270 -300
rect 290 -280 330 -270
rect 290 -300 300 -280
rect 320 -300 330 -280
rect 290 -310 330 -300
<< viali >>
rect 130 420 150 495
rect -25 30 -5 50
rect 145 30 165 50
rect -45 -300 -25 -280
rect 300 -300 320 -280
<< metal1 >>
rect -95 495 330 505
rect -95 420 130 495
rect 150 420 330 495
rect -95 410 330 420
rect -95 50 330 70
rect -95 30 -25 50
rect -5 30 145 50
rect 165 30 330 50
rect -95 10 330 30
rect -95 -280 330 -220
rect -95 -300 -45 -280
rect -25 -300 300 -280
rect 320 -300 330 -280
rect -95 -315 330 -300
<< labels >>
rlabel metal1 -95 40 -95 40 7 clk
port 6 w
rlabel metal1 -95 -270 -95 -270 7 VN
port 7 w
rlabel locali 330 515 330 515 3 Q
port 3 e
rlabel metal1 -95 455 -95 455 7 VP
port 1 w
rlabel locali -95 515 -95 515 7 D
port 2 w
rlabel locali 330 180 330 180 3 QBar
port 4 e
rlabel locali -95 180 -95 180 7 DBar
port 5 w
<< end >>
