magic
tech sky130A
timestamp 1758595984
<< nwell >>
rect -115 -200 155 -60
<< nmos >>
rect 5 -335 20 -235
rect 70 -335 85 -235
<< pmos >>
rect 5 -180 20 -80
rect 70 -180 85 -80
<< ndiff >>
rect -45 -250 5 -235
rect -45 -320 -30 -250
rect -10 -320 5 -250
rect -45 -335 5 -320
rect 20 -335 70 -235
rect 85 -250 135 -235
rect 85 -320 100 -250
rect 120 -320 135 -250
rect 85 -335 135 -320
<< pdiff >>
rect -45 -95 5 -80
rect -45 -165 -30 -95
rect -10 -165 5 -95
rect -45 -180 5 -165
rect 20 -95 70 -80
rect 20 -165 35 -95
rect 55 -165 70 -95
rect 20 -180 70 -165
rect 85 -95 135 -80
rect 85 -165 100 -95
rect 120 -165 135 -95
rect 85 -180 135 -165
<< ndiffc >>
rect -30 -320 -10 -250
rect 100 -320 120 -250
<< pdiffc >>
rect -30 -165 -10 -95
rect 35 -165 55 -95
rect 100 -165 120 -95
<< psubdiff >>
rect -95 -250 -45 -235
rect -95 -320 -80 -250
rect -60 -320 -45 -250
rect -95 -335 -45 -320
<< nsubdiff >>
rect -95 -95 -45 -80
rect -95 -165 -80 -95
rect -60 -165 -45 -95
rect -95 -180 -45 -165
<< psubdiffcont >>
rect -80 -320 -60 -250
<< nsubdiffcont >>
rect -80 -165 -60 -95
<< poly >>
rect 5 -80 20 -65
rect 70 -80 85 -65
rect 5 -235 20 -180
rect 70 -235 85 -180
rect 5 -350 20 -335
rect 70 -350 85 -335
rect -20 -360 20 -350
rect -20 -380 -10 -360
rect 10 -380 20 -360
rect -20 -390 20 -380
rect 45 -360 85 -350
rect 45 -380 55 -360
rect 75 -380 85 -360
rect 45 -390 85 -380
<< polycont >>
rect -10 -380 10 -360
rect 55 -380 75 -360
<< locali >>
rect -90 -95 0 -85
rect -90 -165 -80 -95
rect -60 -165 -30 -95
rect -10 -165 0 -95
rect -90 -175 0 -165
rect 25 -95 65 -85
rect 25 -165 35 -95
rect 55 -165 65 -95
rect 25 -195 65 -165
rect 90 -95 130 -85
rect 90 -165 100 -95
rect 120 -165 130 -95
rect 90 -175 130 -165
rect 25 -220 130 -195
rect -90 -250 0 -240
rect -90 -320 -80 -250
rect -60 -320 -30 -250
rect -10 -320 0 -250
rect -90 -330 0 -320
rect 90 -250 130 -220
rect 90 -320 100 -250
rect 120 -320 130 -250
rect 90 -330 130 -320
rect -20 -360 20 -350
rect -20 -370 -10 -360
rect -115 -380 -10 -370
rect 10 -380 20 -360
rect -115 -390 20 -380
rect 45 -360 85 -350
rect 45 -380 55 -360
rect 75 -380 85 -360
rect 45 -390 85 -380
rect 110 -370 130 -330
rect 110 -390 155 -370
rect 65 -410 85 -390
rect -115 -430 85 -410
<< viali >>
rect -80 -165 -60 -95
rect -30 -165 -10 -95
rect 100 -165 120 -95
rect -80 -320 -60 -250
rect -30 -320 -10 -250
<< metal1 >>
rect -115 -95 155 -85
rect -115 -165 -80 -95
rect -60 -165 -30 -95
rect -10 -165 100 -95
rect 120 -165 155 -95
rect -115 -175 155 -165
rect -115 -250 155 -240
rect -115 -320 -80 -250
rect -60 -320 -30 -250
rect -10 -320 155 -250
rect -115 -330 155 -320
<< labels >>
rlabel locali -115 -420 -115 -420 7 A
port 2 w
rlabel locali -115 -380 -115 -380 7 B
port 3 w
rlabel locali 155 -380 155 -380 3 Y
port 4 e
rlabel metal1 -115 -130 -115 -130 7 VP
port 1 w
rlabel metal1 -115 -285 -115 -285 7 VN
port 5 w
<< end >>
