magic
tech sky130A
timestamp 1758596537
<< nwell >>
rect -195 195 10 335
<< nmos >>
rect -75 60 -60 160
<< pmos >>
rect -75 215 -60 315
<< ndiff >>
rect -125 145 -75 160
rect -125 75 -110 145
rect -90 75 -75 145
rect -125 60 -75 75
rect -60 145 -10 160
rect -60 75 -45 145
rect -25 75 -10 145
rect -60 60 -10 75
<< pdiff >>
rect -125 300 -75 315
rect -125 230 -110 300
rect -90 230 -75 300
rect -125 215 -75 230
rect -60 300 -10 315
rect -60 230 -45 300
rect -25 230 -10 300
rect -60 215 -10 230
<< ndiffc >>
rect -110 75 -90 145
rect -45 75 -25 145
<< pdiffc >>
rect -110 230 -90 300
rect -45 230 -25 300
<< psubdiff >>
rect -175 145 -125 160
rect -175 75 -160 145
rect -140 75 -125 145
rect -175 60 -125 75
<< nsubdiff >>
rect -175 300 -125 315
rect -175 230 -160 300
rect -140 230 -125 300
rect -175 215 -125 230
<< psubdiffcont >>
rect -160 75 -140 145
<< nsubdiffcont >>
rect -160 230 -140 300
<< poly >>
rect -75 315 -60 330
rect -75 160 -60 215
rect -75 45 -60 60
rect -100 35 -60 45
rect -100 15 -90 35
rect -70 15 -60 35
rect -100 5 -60 15
<< polycont >>
rect -90 15 -70 35
<< locali >>
rect -170 300 -80 310
rect -170 230 -160 300
rect -140 230 -110 300
rect -90 230 -80 300
rect -170 220 -80 230
rect -55 300 -15 310
rect -55 230 -45 300
rect -25 230 -15 300
rect -55 220 -15 230
rect -35 155 -15 220
rect -170 145 -80 155
rect -170 75 -160 145
rect -140 75 -110 145
rect -90 75 -80 145
rect -170 65 -80 75
rect -55 145 -15 155
rect -55 75 -45 145
rect -25 75 -15 145
rect -55 65 -15 75
rect -100 35 -60 45
rect -100 25 -90 35
rect -195 15 -90 25
rect -70 15 -60 35
rect -195 5 -60 15
rect -35 25 -15 65
rect -35 5 10 25
<< viali >>
rect -160 230 -140 300
rect -110 230 -90 300
rect -160 75 -140 145
rect -110 75 -90 145
<< metal1 >>
rect -195 300 10 310
rect -195 230 -160 300
rect -140 230 -110 300
rect -90 230 10 300
rect -195 220 10 230
rect -195 145 10 155
rect -195 75 -160 145
rect -140 75 -110 145
rect -90 75 10 145
rect -195 65 10 75
<< labels >>
rlabel locali -195 15 -195 15 7 A
port 2 w
rlabel locali 10 15 10 15 3 Y
port 3 e
rlabel metal1 -195 265 -195 265 7 VP
port 1 w
rlabel metal1 -195 110 -195 110 7 VN
port 4 w
<< end >>
